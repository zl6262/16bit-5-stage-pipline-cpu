`include"define.v"
module reg_data_led(
		input wire sel,
		input wire reg_sel,
		output wire reg_data
);


endmodule 